module ALU(A, B, F, ALU_OP, ZF, OF);
  input [31:0] A, B;       // 输入操作数 A 和 B，每个操作数为 32 位
  input [2:0] ALU_OP;      // 输入 ALU 操作码，用于选择执行的操作
  output reg ZF, OF;       // 输出零标志位 ZF 和溢出标志位 OF
  output reg [31:0] F;     // 输出结果 F，为 32 位

  reg C32;                // 进位标志位 C32

  always @(*) begin       // 组合逻辑块，根据输入信号执行相应操作
    OF = 1'b0;            // 初始化溢出标志位为 0
    C32 = 1'b0;           // 初始化进位标志位为 0

    case (ALU_OP)         // 根据 ALU 操作码选择执行的操作
      3'b000: F = A & B;                  // 操作码为 000，执行 A 与 B 的按位与操作
      3'b001: F = A | B;                  // 操作码为 001，执行 A 与 B 的按位或操作
      3'b010: F = A ^ B;                  // 操作码为 010，执行 A 与 B 的按位异或操作
      3'b011: F = ~(A ^ B);               // 操作码为 011，执行 A 与 B 的按位异或后取反操作
      3'b100: begin                       // 操作码为 100，执行 A 与 B 的加法操作
        {C32, F} = A + B;                 // 将 A 和 B 相加，进位结果存储在 C32，和存储在 F
        OF = A[31] ^ B[31] ^ F[31] ^ C32;  // 计算溢出标志位 OF
      end
      3'b101: begin                       // 操作码为 101，执行 A 与 B 的减法操作
        {C32, F} = A - B;                 // 将 A 减去 B，进位结果存储在 C32，差存储在 F
        OF = A[31] ^ B[31] ^ F[31] ^ C32;  // 计算溢出标志位 OF
      end
      3'b110:                            // 操作码为 110，执行 A 与 B 的比较操作
        if (A < B)                       // 如果 A 小于 B
          F = 1;                         // 将结果 F 设置为 1
        else
          F = 0;                         // 否则将结果 F 设置为 0
      3'b111: F = B << A;                 // 操作码为 111，执行 B 的左移 A 位操作
    endcase

    if (F == 0)
      ZF = 1;                           // 如果结果 F 等于 0，将零标志位 ZF 设置为 1
    else
      ZF = 0;                           // 否则将零标志位 ZF 设置为 0
  end
endmodule
